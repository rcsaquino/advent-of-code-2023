module day_01

pub fn print_answers(input string) {
	println("---DAY 1---")
	println("Part 1: ${part_one(input)}")
	println("Part 2: ${part_two(input)}")
}
