module day_01

pub fn solution(input string) {
	lines := input.split('\r\n')

	println('Part 1: ${part_one(lines)}')
	println('Part 2: ${part_two(lines)}')
}
